-- Random Access Memory with 1 read/write port

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- RAM entity
ENTITY RANDOM_ACCESS_MEMORY IS
  PORT(
    DATAIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    W_R : IN STD_LOGIC; --! Write when 0, Read when 1
    DATAOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END ENTITY;

-- RAM architecture
ARCHITECTURE RAM_BEHAVIOUR OF RANDOM_ACCESS_MEMORY IS

TYPE RAM_MEM IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL MEMORY : RAM_MEM;
SIGNAL ADDR : INTEGER RANGE 0 TO 31;

BEGIN

  PROCESS(ADDRESS, DATAIN, W_R)
  BEGIN
    ADDR<=CONV_INTEGER(ADDRESS);
    IF(W_R='0') THEN
      MEMORY(ADDR)<=DATAIN;
    ELSIF(W_R='1') THEN
      DATAOUT<=MEMORY(ADDR);
    ELSE
      DATAOUT<="00000000000000000000000000000000";
    END IF;
  END PROCESS;

END RAM_BEHAVIOR;
